`default_nettype none

module vga_image(
    input wire clk_in,
    input wire reset,
    output reg r1,
    output reg r2,
    output reg b1,
    output reg b2,
    output reg g1,
    output reg g2,
    output wire h_sync,
    output wire v_sync,
    output wire led,
    output wire locked_led
  );

wire clk_sys;
wire display_en;
//reg [9:0] h_count;
wire [9:0] h_count;
//reg [9:0] v_count;
wire [9:0] v_count;
assign  led = clk_sys;


// RAM interfacing
// 510 x 85
localparam  AddressWidth = 9; // 2^7 = 128
localparam  DataWidth = 512;
reg [AddressWidth-1:0] addr;
reg [AddressWidth-1:0] addr_counter = 0;
reg [DataWidth-1:0]  data_in;
reg [DataWidth-1:0]  data_out;

reg [DataWidth-1:0]  pixel_row_current;
reg [DataWidth-1:0]  pixel_row_next;

reg [6-1:0]  rgb_out = 5'h3F;

reg rw = 1; // Set enabled read of RAM


localparam  h_total  = 480;
localparam  v_total  = 640;
localparam  h_image_pixel = 85;
localparam  v_image_pixel = 116;

localparam   h_image_start = 198;
localparam   h_image_finish = 283;
localparam   v_image_start = 262;
localparam   v_image_finish = 378;

// Draw in the frame the image, canvas otherwise
always @(posedge clk_sys) begin
  if (display_en) begin
      if ((v_count > v_image_start-1 && v_count < v_image_finish-1)
       && (h_count > h_image_start-1 && h_count < h_image_finish-1))
        begin
        //Image
        r1 <= rgb_out[0];
        r2 <= rgb_out[1];
        g1 <= rgb_out[2];
        g2 <= rgb_out[3];
        b1 <= rgb_out[4];
        b2 <= rgb_out[5];
        /*
        r1 <= 1'b1;
        r2 <= 1'b1;
        g1 <= 1'b1;
        g2 <= 1'b1;
        b1 <= 1'b0;
        b2 <= 1'b0;
        */
        end
    else begin
      //Canvas color
      r1 <= 1'b1;
      r2 <= 1'b0;
      g1 <= 1'b1;
      g2 <= 1'b0;
      b1 <= 1'b1;
      b2 <= 1'b1;
    end
  end
  else begin
  // Pixels out of display
  r1 <= 1'b0;
  r2 <= 1'b0;
  g1 <= 1'b0;
  g2 <= 1'b0;
  b1 <= 1'b0;
  b2 <= 1'b0;
  end
end

/*
always @(clk_sys)begin
  if (reset)
    addr_counter <= 0;
  else begin
    if (v_counter > v_image_start-1 && (h_counter > h_image_start && h_counter < h_image_finish))
    if (addr_counter >= 116)
      addr_counter <= 0;
    else
      addr_counter <= addr_counter + 1;
    end
end
*/


vga_sync vga_s(
      .clk_in(clk_in),         //12MHz clock input
      .reset(reset),           // RST assigned to SW1
      .h_sync(h_sync),
      .v_sync(v_sync),
      .clk_sys(clk_sys),       //25.125 MHz clock generated by PLL
      .h_count(h_count),
      .v_count(v_count),
      .display_en(display_en), // '1' => pixel region
      .locked(locked_led)      // PLL signal, '1' => OK
      );


ram #(
       .AddressWidth(AddressWidth),
       .DataWidth(DataWidth)
      )ram
      (
       .clk(clk_sys),
       .rw(rw), //Read '1', write '0'
       .addr(addr),
       .data_in(data_in),
       .data_out(data_out)
       );


endmodule
