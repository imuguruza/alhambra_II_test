// Copyright 2020 Iñigo Muguruza Goenaga
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

/*
  VGA IMAGE module
  ================

  - Instantiates vga_sync for sync signal generation
  - Creates canvas color
  - Reads RAM memory and displays image in pixel range
  - Lokecd Led => Shows if PLL is working right, debugging purposes
  - CLK LED => LED assigned to 25MHz clock, debugging purposes
  - Color format: RRRGGBB

*/
`default_nettype none

module vga_image(
    input wire clk_in,
    input wire reset,
    output reg [8:0] rgb_port,
    output wire h_sync,
    output wire v_sync,
    output wire clk_led,
    output wire locked_led
  );

wire clk_sys;
wire display_en;
//reg [9:0] h_count;
wire [9:0] h_count;
//reg [9:0] v_count;
wire [9:0] v_count;


// RAM interfacing
// (100 pixel x 8 bits color) x 100 pixel
localparam  AddressWidth = 14; // 2^14 = 16384
localparam  DataWidth = 8; //
reg [AddressWidth-1:0] addr = 0;
reg [DataWidth-1:0]  data_in;
//reg [DataWidth-1:0]  data_out;
wire [DataWidth-1:0]  w_data_out;

reg [7:0]  rgb_out;

reg rw = 1; // Set enabled read of RAM


localparam  h_total  = 640;
localparam  v_total  = 480;
localparam  h_image_pixel = 100;
localparam  v_image_pixel = 100;

localparam addr_amount = 10000; // Total pixel amount 100x100

// Calculate where the image nees to be drawn
localparam   h_image_start = h_total/2 - h_image_pixel/2;
localparam   h_image_finish = h_total/2 + h_image_pixel/2;
localparam   v_image_start = v_total/2 - v_image_pixel/2;
localparam   v_image_finish = v_total/2 + v_image_pixel/2;

// Load the image from RAM
always @(posedge clk_sys) begin
      if ((v_count >= v_image_start-1 && v_count < v_image_finish-1)
       && (h_count >= h_image_start-1 && h_count < h_image_finish-1))
       begin
        //Load Image from RAM
        rgb_out <= w_data_out;
        addr <= addr + 1;//Load new row pixel
        if (addr >= addr_amount -1)//Out of bounce, go to 0
          addr <= 0;
      end
end

// Draw in the frame the image, canvas otherwise
always @(posedge clk_sys) begin
  if (display_en) begin
      if ((v_count > v_image_start-1 && v_count < v_image_finish-1)
       && (h_count > h_image_start-1 && h_count < h_image_finish-1))
        //Image
        rgb_port <= {1'b1,rgb_out};
      else
      rgb_port <= 9'b10111111;
  end else
  // Pixels out of display
  rgb_port <= 9'b000000000;
end


//Blink Led with clk
assign  clk_led = clk_sys;

vga_sync vga_s(
      .clk_in(clk_in),         //12MHz clock input
      .reset(reset),           // RST assigned to SW1
      .h_sync(h_sync),
      .v_sync(v_sync),
      .clk_sys(clk_sys),       //25.125 MHz clock generated by PLL
      .h_count(h_count),
      .v_count(v_count),
      .display_en(display_en), // '1' => pixel region
      .locked(locked_led)      // PLL signal, '1' => OK
      );

ram #(
       .AddressWidth(AddressWidth),
       .DataWidth(DataWidth),
       .RAMFILE("bender.mem")
      )ram
      (
       .clk(clk_sys),
       .rw(rw), //Read '1', write '0'
       .addr(addr),
       .data_in(data_in),
       .data_out(w_data_out)
       );


endmodule
