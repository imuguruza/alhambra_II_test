// Hz
`define F_100Hz   120_000
`define F_50Hz   240_000
`define F_40Hz   300_000
`define F_20Hz   600_000
`define F_10Hz   1_200_000
`define F_8Hz   1_500_000
`define F_4Hz   3_000_000
`define F_2Hz   6_000_000
`define F_1Hz   12_000_000
